CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
490 0 1 200 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
10
9 CC 7-Seg~
183 962 77 0 18 19
10 10 9 8 7 6 5 4 17 18
1 1 1 0 0 1 1 2 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5130 0 0
2
5.89883e-315 0
0
6 74LS48
188 794 197 0 14 29
0 11 13 12 2 19 20 4 5 6
7 8 9 10 21
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
391 0 0
2
5.89883e-315 5.26354e-315
0
9 2-In AND~
219 630 146 0 3 22
0 14 13 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3124 0 0
2
5.89883e-315 5.30499e-315
0
9 2-In AND~
219 484 137 0 3 22
0 2 12 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3421 0 0
2
5.89883e-315 5.32571e-315
0
2 +V
167 261 187 0 1 3
0 3
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
5.89883e-315 5.34643e-315
0
7 Pulser~
4 164 321 0 10 12
0 22 23 24 15 0 0 5 5 4
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5572 0 0
2
43530.3 0
0
6 74112~
219 697 277 0 7 32
0 3 16 15 16 3 25 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8901 0 0
2
43530.3 1
0
6 74112~
219 549 277 0 7 32
0 3 14 15 14 3 26 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7361 0 0
2
43530.3 2
0
6 74112~
219 394 303 0 7 32
0 3 2 15 2 3 27 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
4747 0 0
2
43530.3 3
0
6 74112~
219 262 300 0 7 32
0 3 28 15 29 3 30 2
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
972 0 0
2
43530.3 4
0
42
2 0 2 0 0 4096 0 9 0 0 10 3
370 267
370 250
360 250
0 0 3 0 0 4096 0 0 0 20 7 2
612 196
612 365
0 0 3 0 0 0 0 0 0 20 7 2
472 196
472 365
0 0 3 0 0 0 0 0 0 20 7 2
315 196
315 365
5 0 3 0 0 0 0 8 0 0 7 2
549 289
549 365
5 0 3 0 0 0 0 9 0 0 7 4
394 315
394 360
395 360
395 365
5 5 3 0 0 8192 0 10 7 0 0 4
262 312
262 365
697 365
697 289
0 4 2 0 0 8320 0 0 2 9 0 3
335 264
335 188
762 188
7 0 2 0 0 0 0 10 0 0 10 2
286 264
360 264
4 1 2 0 0 0 0 9 4 0 0 4
370 285
360 285
360 128
460 128
7 0 4 0 0 4096 0 1 0 0 27 2
977 113
978 113
6 0 5 0 0 4096 0 1 0 0 28 2
971 113
972 113
5 0 6 0 0 4096 0 1 0 0 29 2
965 113
966 113
4 0 7 0 0 4096 0 1 0 0 30 2
959 113
960 113
3 0 8 0 0 4096 0 1 0 0 31 2
953 113
954 113
2 0 9 0 0 4096 0 1 0 0 32 2
947 113
948 113
1 0 10 0 0 4096 0 1 0 0 33 2
941 113
942 113
1 0 3 0 0 0 0 8 0 0 20 2
549 214
549 196
1 0 3 0 0 0 0 9 0 0 20 2
394 240
394 196
1 1 3 0 0 4224 0 5 7 0 0 3
261 196
697 196
697 214
1 1 3 0 0 0 0 10 5 0 0 3
262 237
261 237
261 196
7 1 11 0 0 8320 0 7 2 0 0 4
721 241
753 241
753 161
762 161
0 3 12 0 0 12416 0 0 2 39 0 4
439 240
458 240
458 179
762 179
0 2 13 0 0 12416 0 0 2 38 0 4
590 241
621 241
621 170
762 170
2 0 14 0 0 4096 0 8 0 0 26 2
525 241
505 241
4 3 14 0 0 8320 0 8 4 0 0 3
525 259
505 259
505 137
7 0 4 0 0 4224 0 2 0 0 0 4
826 161
978 161
978 110
979 110
8 0 5 0 0 4224 0 2 0 0 0 4
826 170
972 170
972 110
973 110
9 0 6 0 0 4224 0 2 0 0 0 4
826 179
966 179
966 110
967 110
10 0 7 0 0 4224 0 2 0 0 0 4
826 188
960 188
960 110
961 110
11 0 8 0 0 4224 0 2 0 0 0 4
826 197
954 197
954 110
955 110
12 0 9 0 0 4224 0 2 0 0 0 4
826 206
948 206
948 110
949 110
13 0 10 0 0 4224 0 2 0 0 0 4
826 215
942 215
942 110
943 110
3 0 15 0 0 8192 0 10 0 0 42 3
232 273
206 273
206 321
3 1 14 0 0 0 0 4 3 0 0 2
505 137
606 137
2 0 16 0 0 4096 0 7 0 0 37 2
673 241
653 241
3 4 16 0 0 8320 0 3 7 0 0 4
651 146
653 146
653 259
673 259
7 2 13 0 0 0 0 8 3 0 0 4
573 241
590 241
590 155
606 155
2 7 12 0 0 0 0 4 9 0 0 4
460 146
439 146
439 267
418 267
3 0 15 0 0 8192 0 8 0 0 42 3
519 250
487 250
487 321
3 0 15 0 0 0 0 9 0 0 42 3
364 276
340 276
340 321
4 3 15 0 0 4224 0 6 7 0 0 4
194 321
641 321
641 250
667 250
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
358 402 553 424
367 410 543 426
22 BOYBOY, JUVENAR JR. C.
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
